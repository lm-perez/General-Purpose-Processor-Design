LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY decod IS
	PORT( w		:IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
				y		:BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0));
END decod;

ARCHITECTURE BEHAVIOR OF decod IS
	SIGNAL Ew: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	Ew <= w;
	WITH Ew SELECT
		y<= "0000000000000001" WHEN "0000",
		"0000000000000010" WHEN "0001",
		"0000000000000100" WHEN "0010",
		"0000000000001000" WHEN "0011",
		"0000000000010000" WHEN "0100",
		"0000000000100000" WHEN "0101",
		"0000000001000000" WHEN "0110",
		"0000000010000000" WHEN "0111",
		"0000000100000000" WHEN "1000",
		
		"0000000000000000" WHEN OTHERS;
				
				
END BEHAVIOR;
